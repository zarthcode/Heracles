
module AbsoluteEncoder ( ADCValue, clk);
	
	
endmodule