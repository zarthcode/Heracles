// Quadature encoder implementation.

module QuadatureEncoder