
module AbsoluteEncoder ( ADCValue, 