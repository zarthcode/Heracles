// Wishbone EFB Master

module efb_master();
	
	
	
	
endmodule