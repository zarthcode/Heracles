// Heracles Device

module Heracles();
	
	// Oscillator
	
		// Clock
		// Trimdac clk
		// spi clk
		// stepper clock
		// servo clk
		
	// I2C Interface
	
	// Config Registers
	
	// SPI Slave Interface
	
	// TrimDAC SPI Bus
	
	// Encoder Channels
	
	// Stepper Channels
	
	// Servo Channels
	
	// PID Channels
	
	
endmodule