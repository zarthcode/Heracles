// Open-loop stepper motor with microstep morphing.

module SmoothStepper();
	
	// Inputs
	
	// Outputs
	
	// Registers
	
	
	
endmodule;